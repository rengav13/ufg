module sensorDePresenca(sinal,led);

input sinal;
output led;
wire led;

assign led=sinal;

endmodule
