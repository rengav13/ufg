library verilog;
use verilog.vl_types.all;
entity teste_GSM_vlg_vec_tst is
end teste_GSM_vlg_vec_tst;
