library verilog;
use verilog.vl_types.all;
entity teste_Mod_comm_vlg_vec_tst is
end teste_Mod_comm_vlg_vec_tst;
